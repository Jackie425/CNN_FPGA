`timescale 1ns / 1ps

module FeatureMapMemoryTop # (

)
(
    
);


endmodule