`timescale 1ns / 1ps

module FeatureMapDRM #(

)
(
    

);



endmodule