`timescale 1ns / 1ps

module FeatureMapCtrl # (
             
)
(
     
);


endmodule
