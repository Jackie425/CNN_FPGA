`timescale 1ns / 1ps

module PWConvPreProcess # (

)
(

);


endmodule